/*
  Eric Villasenor
  evillase@gmail.com

  register file test bench
*/

// mapped needs this
`include "register_file_if.vh"

// mapped timing needs this. 1ns is too fast
`timescale 1 ns / 1 ns

module register_file_tb;

  parameter PERIOD = 10;

  logic CLK = 0, nRST;

  // test vars
  int v1 = 1;
  int v2 = 4721;
  int v3 = 25119;

  // clock
  always #(PERIOD/2) CLK++;

  // interface
  register_file_if rfif ();//
  // test program
   test PROG (.CLK(CLK), .nRST(nRST), .rfif(rfif));   

   
  // DUT
`ifndef MAPPED
  register_file DUT(CLK, nRST, rfif);
`else
  register_file DUT(
    .\rfif.rdat2 (rfif.rdat2),
    .\rfif.rdat1 (rfif.rdat1),
    .\rfif.wdat (rfif.wdat),
    .\rfif.rsel2 (rfif.rsel2),
    .\rfif.rsel1 (rfif.rsel1),
    .\rfif.wsel (rfif.wsel),
    .\rfif.WEN (rfif.WEN),
    .\nRST (nRST),
    .\CLK (CLK)
  );
`endif

endmodule

program test
import cpu_types_pkg::*;
(
   input logic CLK,
   output logic nRST,
   register_file_if.tb rfif
 );

 parameter PERIOD=10;

initial 
begin
 
   word_t data_in [32];
   
 
   data_in[0]='0;
   nRST=0;
   #(PERIOD/2);      
   rfif.wdat='0;
   rfif.rsel1='0;
   rfif.rsel2='0;
   rfif.wsel='0;
   rfif.WEN=0;
   nRST=1;
   #(PERIOD);
   
   /////////////////////////////
   rfif.wdat=123;
   rfif.rsel1=0;
   rfif.rsel2=0;
   rfif.wsel=1;
   rfif.WEN=1;
   #(PERIOD);
   
      $display("rdat1 and rdat2 value");
   assert(rfif.rdat1==0 && rfif.rdat2 ==0)
     else begin
	$error("case 1 wrong");
     end
////////////////////////// write to 1 and load from 1 /////////////////            

      rfif.wdat=4567;
      rfif.rsel1=1;
      rfif.rsel2=1;
      rfif.wsel=2;
      rfif.WEN=1;
      #(PERIOD);
     assert(rfif.rdat1==123 && rfif.rdat2 ==123)
     $display("write to 2 and read from 1");
     else begin
	$error("case 2 wrong : write to 2 and reading from 1");
     end
///////////////// write to 2 and load from 1 and 2 ///////////////////

      
 
      rfif.wdat=19949;
      rfif.rsel1=1;
      rfif.rsel2=2;
      rfif.wsel=31;
      rfif.WEN=1;
      #(PERIOD);
      $display("write/read from 1 and 2");
     assert(rfif.rdat1==123 && rfif.rdat2 ==4567)
     else begin
	$error("case 3 wrong : writing/reading from 1 and 2");
     end
///////////////////// don't write, just read/////////////////////////////   
      rfif.wdat=0;
      rfif.rsel1=2;
      rfif.rsel2=31;
      rfif.wsel=0;
      rfif.WEN=0;
      #(PERIOD);
     assert(rfif.rdat1==4567 && rfif.rdat2 ==19949)
     else begin
	$error("case 4 wrong : no write / reading from 30 and 31");
     end
//////////////////////////////////////////////////////////////////
      rfif.wdat=9876;
      rfif.rsel1=0;
      rfif.rsel2=0;
      rfif.wsel=0;
      rfif.WEN=1;
      #(PERIOD);
      rfif.wdat=0;
      rfif.rsel1=0;
      rfif.rsel2=0;
      rfif.wsel=0;
      rfif.WEN=0;
   #(PERIOD);   
   
end
   
//       
endprogram
